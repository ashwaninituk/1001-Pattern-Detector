magic
tech scmos
timestamp 1606150958
<< nwell >>
rect -98 26 307 72
<< polysilicon >>
rect -92 63 -90 74
rect -84 63 -82 65
rect -76 63 -74 74
rect -68 63 -66 65
rect -60 63 -58 74
rect -52 63 -50 65
rect -34 51 -32 53
rect -26 51 -24 88
rect -18 51 -16 81
rect -10 51 -8 53
rect 25 51 27 53
rect 33 51 35 81
rect 41 51 43 88
rect 49 51 51 53
rect 5 39 7 41
rect 83 49 85 74
rect 109 51 111 74
rect 117 51 119 53
rect 134 51 136 53
rect 142 51 144 88
rect 150 51 152 81
rect 158 51 160 53
rect 193 51 195 53
rect 201 51 203 81
rect 209 51 211 88
rect 217 51 219 53
rect 63 39 65 41
rect 101 39 103 41
rect 173 39 175 41
rect 251 49 253 74
rect 267 63 269 74
rect 275 63 277 65
rect 283 63 285 74
rect 231 39 233 41
rect 299 39 301 41
rect -92 12 -90 27
rect -84 12 -82 27
rect -76 12 -74 27
rect -68 12 -66 27
rect -60 12 -58 27
rect -52 12 -50 27
rect -34 22 -32 27
rect -26 25 -24 27
rect -18 25 -16 27
rect -34 12 -32 18
rect -10 17 -8 27
rect 5 24 7 27
rect -26 12 -24 14
rect -18 12 -16 14
rect -10 12 -8 13
rect 5 12 7 20
rect 25 17 27 27
rect 33 25 35 27
rect 41 25 43 27
rect 49 17 51 27
rect 63 24 65 27
rect 83 25 85 27
rect 25 12 27 13
rect 33 12 35 14
rect 41 12 43 14
rect 49 12 51 13
rect 63 12 65 20
rect 101 12 103 27
rect 109 12 111 27
rect 117 12 119 27
rect 134 25 136 27
rect 142 25 144 27
rect 150 25 152 27
rect 134 12 136 21
rect 158 17 160 27
rect 173 24 175 27
rect 142 12 144 14
rect 150 12 152 14
rect 158 12 160 13
rect 173 12 175 20
rect 193 17 195 27
rect 201 25 203 27
rect 209 25 211 27
rect 217 17 219 27
rect 231 24 233 27
rect 251 25 253 27
rect 193 12 195 13
rect 201 12 203 14
rect 209 12 211 14
rect 217 12 219 13
rect 231 12 233 20
rect 267 12 269 27
rect 275 12 277 27
rect 283 12 285 27
rect 299 19 301 27
rect 300 15 301 19
rect 299 12 301 15
rect 5 4 7 6
rect 63 4 65 6
rect 173 4 175 6
rect 231 4 233 6
rect 267 4 269 6
rect -92 -2 -90 0
rect -84 -11 -82 0
rect -76 -2 -74 0
rect -68 -11 -66 0
rect -60 -2 -58 0
rect -52 -11 -50 0
rect -34 -2 -32 0
rect -26 -18 -24 0
rect -18 -25 -16 0
rect -10 -2 -8 0
rect 25 -2 27 0
rect 33 -25 35 0
rect 41 -18 43 0
rect 49 -2 51 0
rect 101 -11 103 0
rect 109 -2 111 0
rect 117 -11 119 0
rect 134 -2 136 0
rect 142 -18 144 0
rect 150 -25 152 0
rect 158 -2 160 0
rect 193 -2 195 0
rect 201 -25 203 0
rect 209 -18 211 0
rect 217 -2 219 0
rect 275 -11 277 6
rect 283 4 285 6
rect 299 4 301 6
<< ndiffusion >>
rect -97 4 -92 12
rect -93 0 -92 4
rect -90 8 -89 12
rect -85 8 -84 12
rect -90 0 -84 8
rect -82 4 -76 12
rect -82 0 -81 4
rect -77 0 -76 4
rect -74 8 -73 12
rect -69 8 -68 12
rect -74 5 -68 8
rect -74 1 -73 5
rect -69 1 -68 5
rect -74 0 -68 1
rect -66 8 -65 12
rect -61 8 -60 12
rect -66 0 -60 8
rect -58 5 -52 12
rect -58 1 -57 5
rect -53 1 -52 5
rect -58 0 -52 1
rect -50 8 -49 12
rect -45 8 -44 12
rect -50 0 -44 8
rect -39 5 -34 12
rect -35 1 -34 5
rect -39 0 -34 1
rect -32 0 -26 12
rect -24 8 -23 12
rect -19 8 -18 12
rect -24 0 -18 8
rect -16 0 -10 12
rect -8 6 5 12
rect 7 10 16 12
rect 7 6 10 10
rect 14 6 16 10
rect -8 5 -1 6
rect -8 1 -7 5
rect -3 1 -1 5
rect 20 5 25 12
rect -8 0 -1 1
rect 24 1 25 5
rect 20 0 25 1
rect 27 0 33 12
rect 35 8 36 12
rect 40 8 41 12
rect 35 0 41 8
rect 43 0 49 12
rect 51 6 63 12
rect 65 10 74 12
rect 65 6 68 10
rect 72 6 74 10
rect 51 5 58 6
rect 51 1 52 5
rect 56 1 58 5
rect 96 4 101 12
rect 51 0 58 1
rect 100 0 101 4
rect 103 6 109 12
rect 103 2 104 6
rect 108 2 109 6
rect 103 0 109 2
rect 111 8 112 12
rect 116 8 117 12
rect 111 0 117 8
rect 119 6 124 12
rect 119 2 120 6
rect 119 0 124 2
rect 129 5 134 12
rect 133 1 134 5
rect 129 0 134 1
rect 136 0 142 12
rect 144 8 145 12
rect 149 8 150 12
rect 144 0 150 8
rect 152 0 158 12
rect 160 6 173 12
rect 175 10 184 12
rect 175 6 178 10
rect 182 6 184 10
rect 160 5 167 6
rect 160 1 161 5
rect 165 1 167 5
rect 188 5 193 12
rect 160 0 167 1
rect 192 1 193 5
rect 188 0 193 1
rect 195 0 201 12
rect 203 8 204 12
rect 208 8 209 12
rect 203 0 209 8
rect 211 0 217 12
rect 219 6 231 12
rect 233 10 242 12
rect 233 6 236 10
rect 240 6 242 10
rect 262 10 267 12
rect 266 6 267 10
rect 269 8 270 12
rect 274 8 275 12
rect 269 6 275 8
rect 277 10 283 12
rect 277 6 278 10
rect 282 6 283 10
rect 285 8 286 12
rect 285 6 290 8
rect 294 10 299 12
rect 298 6 299 10
rect 301 8 302 12
rect 301 6 306 8
rect 219 5 226 6
rect 219 1 220 5
rect 224 1 226 5
rect 219 0 226 1
<< pdiffusion >>
rect -93 59 -92 63
rect -97 27 -92 59
rect -90 27 -84 63
rect -82 27 -76 63
rect -74 31 -68 63
rect -74 27 -73 31
rect -69 27 -68 31
rect -66 27 -60 63
rect -58 27 -52 63
rect -50 59 -49 63
rect -45 59 -44 63
rect -50 27 -44 59
rect -39 49 -34 51
rect -35 45 -34 49
rect -39 27 -34 45
rect -32 27 -26 51
rect -24 33 -18 51
rect -24 29 -23 33
rect -19 29 -18 33
rect -24 27 -18 29
rect -16 27 -10 51
rect -8 49 -1 51
rect -8 45 -7 49
rect -3 45 -1 49
rect -8 39 -1 45
rect 20 49 25 51
rect 24 45 25 49
rect -8 27 5 39
rect 7 31 16 39
rect 7 27 10 31
rect 14 27 16 31
rect 20 27 25 45
rect 27 27 33 51
rect 35 33 41 51
rect 35 29 36 33
rect 40 29 41 33
rect 35 27 41 29
rect 43 27 49 51
rect 51 49 58 51
rect 51 45 52 49
rect 56 45 58 49
rect 51 39 58 45
rect 78 43 83 49
rect 82 39 83 43
rect 51 27 63 39
rect 65 31 74 39
rect 65 27 68 31
rect 72 27 74 31
rect 78 27 83 39
rect 85 45 86 49
rect 85 27 90 45
rect 106 39 109 51
rect 100 35 101 39
rect 96 27 101 35
rect 103 31 109 39
rect 103 27 104 31
rect 108 27 109 31
rect 111 27 117 51
rect 119 47 120 51
rect 119 27 124 47
rect 129 49 134 51
rect 133 45 134 49
rect 129 27 134 45
rect 136 27 142 51
rect 144 33 150 51
rect 144 29 145 33
rect 149 29 150 33
rect 144 27 150 29
rect 152 27 158 51
rect 160 49 167 51
rect 160 45 161 49
rect 165 45 167 49
rect 160 39 167 45
rect 188 49 193 51
rect 192 45 193 49
rect 160 27 173 39
rect 175 31 184 39
rect 175 27 178 31
rect 182 27 184 31
rect 188 27 193 45
rect 195 27 201 51
rect 203 33 209 51
rect 203 29 204 33
rect 208 29 209 33
rect 203 27 209 29
rect 211 27 217 51
rect 219 49 226 51
rect 266 59 267 63
rect 219 45 220 49
rect 224 45 226 49
rect 219 39 226 45
rect 246 43 251 49
rect 250 39 251 43
rect 219 27 231 39
rect 233 31 242 39
rect 233 27 236 31
rect 240 27 242 31
rect 246 27 251 39
rect 253 45 254 49
rect 253 27 258 45
rect 262 27 267 59
rect 269 27 275 63
rect 277 27 283 63
rect 285 31 290 63
rect 285 27 286 31
rect 298 35 299 39
rect 294 27 299 35
rect 301 31 306 39
rect 301 27 302 31
<< metal1 >>
rect -112 88 -28 92
rect -24 88 41 92
rect 45 88 140 92
rect 144 88 209 92
rect -112 -25 -109 88
rect -106 81 -18 85
rect -14 81 32 85
rect 36 81 150 85
rect 154 81 199 85
rect -106 -18 -103 81
rect -98 74 -95 78
rect -82 74 -78 78
rect -66 74 -62 78
rect 78 74 81 78
rect 105 74 107 78
rect 246 74 249 78
rect 262 74 265 78
rect 277 74 281 78
rect -93 67 -49 71
rect -45 67 -39 71
rect -35 67 20 71
rect 24 67 86 71
rect 90 67 96 71
rect 100 67 120 71
rect 124 67 129 71
rect 133 67 188 71
rect 192 67 254 71
rect 258 67 262 71
rect 266 67 294 71
rect -97 63 -94 67
rect -48 63 -45 67
rect -39 49 -36 67
rect -7 49 -3 67
rect 20 49 23 67
rect 52 49 56 67
rect 87 49 90 67
rect 58 39 78 42
rect 96 39 99 67
rect 121 51 124 67
rect 129 49 132 67
rect 161 49 165 67
rect 188 49 191 67
rect 220 49 224 67
rect 255 49 258 67
rect 262 63 265 67
rect 226 39 246 42
rect 294 39 298 67
rect -72 22 -69 27
rect -23 24 -20 29
rect -72 19 -36 22
rect -65 12 -62 19
rect -49 18 -36 19
rect -23 20 3 24
rect -49 12 -46 18
rect -23 12 -20 20
rect 10 16 13 27
rect 36 24 39 29
rect 58 24 61 39
rect 36 20 61 24
rect 68 20 71 27
rect 105 25 108 27
rect 105 21 132 25
rect 145 24 148 29
rect -6 13 23 16
rect -85 9 -73 12
rect 10 10 13 13
rect 36 12 39 20
rect 68 16 78 20
rect 53 13 71 16
rect 68 10 71 13
rect 112 12 115 21
rect 145 20 171 24
rect 145 12 148 20
rect 178 16 181 27
rect 204 24 207 29
rect 226 24 229 39
rect 204 20 229 24
rect 236 20 239 27
rect 287 24 290 27
rect 271 21 292 24
rect 162 13 191 16
rect 178 10 181 13
rect 204 12 207 20
rect 236 16 246 20
rect 221 13 239 16
rect 236 10 239 13
rect 271 12 274 21
rect 287 20 292 21
rect 287 12 290 20
rect 303 19 306 27
rect 295 15 296 19
rect 303 15 308 19
rect 303 12 306 15
rect -69 1 -57 4
rect -97 -4 -94 0
rect -81 -4 -78 0
rect -39 -4 -36 1
rect -7 -4 -3 1
rect 20 -4 23 1
rect 52 -4 56 1
rect 108 2 120 5
rect 96 -4 99 0
rect 129 -4 132 1
rect 161 -4 165 1
rect 188 -4 191 1
rect 220 -4 224 1
rect 262 -4 265 6
rect 279 -4 282 6
rect 294 -4 298 6
rect -93 -8 -81 -4
rect -77 -8 -39 -4
rect -35 -8 -7 -4
rect -3 -8 20 -4
rect 24 -8 52 -4
rect 56 -8 96 -4
rect 100 -8 129 -4
rect 133 -8 161 -4
rect 165 -8 188 -4
rect 192 -8 220 -4
rect 224 -8 262 -4
rect 266 -8 294 -4
rect -89 -15 -86 -11
rect -64 -15 -61 -11
rect -48 -15 -45 -11
rect 97 -15 99 -11
rect 113 -15 115 -11
rect 270 -15 273 -11
rect -106 -22 -28 -18
rect -24 -22 40 -18
rect 44 -22 140 -18
rect 144 -22 209 -18
rect -112 -29 -18 -25
rect -14 -29 31 -25
rect 35 -29 150 -25
rect 154 -29 199 -25
<< ntransistor >>
rect -92 0 -90 12
rect -84 0 -82 12
rect -76 0 -74 12
rect -68 0 -66 12
rect -60 0 -58 12
rect -52 0 -50 12
rect -34 0 -32 12
rect -26 0 -24 12
rect -18 0 -16 12
rect -10 0 -8 12
rect 5 6 7 12
rect 25 0 27 12
rect 33 0 35 12
rect 41 0 43 12
rect 49 0 51 12
rect 63 6 65 12
rect 101 0 103 12
rect 109 0 111 12
rect 117 0 119 12
rect 134 0 136 12
rect 142 0 144 12
rect 150 0 152 12
rect 158 0 160 12
rect 173 6 175 12
rect 193 0 195 12
rect 201 0 203 12
rect 209 0 211 12
rect 217 0 219 12
rect 231 6 233 12
rect 267 6 269 12
rect 275 6 277 12
rect 283 6 285 12
rect 299 6 301 12
<< ptransistor >>
rect -92 27 -90 63
rect -84 27 -82 63
rect -76 27 -74 63
rect -68 27 -66 63
rect -60 27 -58 63
rect -52 27 -50 63
rect -34 27 -32 51
rect -26 27 -24 51
rect -18 27 -16 51
rect -10 27 -8 51
rect 5 27 7 39
rect 25 27 27 51
rect 33 27 35 51
rect 41 27 43 51
rect 49 27 51 51
rect 63 27 65 39
rect 83 27 85 49
rect 101 27 103 39
rect 109 27 111 51
rect 117 27 119 51
rect 134 27 136 51
rect 142 27 144 51
rect 150 27 152 51
rect 158 27 160 51
rect 173 27 175 39
rect 193 27 195 51
rect 201 27 203 51
rect 209 27 211 51
rect 217 27 219 51
rect 231 27 233 39
rect 251 27 253 49
rect 267 27 269 63
rect 275 27 277 63
rect 283 27 285 63
rect 299 27 301 39
<< polycontact >>
rect -28 88 -24 92
rect -95 74 -90 78
rect -78 74 -74 78
rect -62 74 -58 78
rect 41 88 45 92
rect 140 88 144 92
rect -18 81 -14 85
rect 32 81 36 85
rect 81 74 85 78
rect 107 74 111 78
rect 209 88 213 92
rect 150 81 154 85
rect 199 81 203 85
rect 249 74 253 78
rect 265 74 269 78
rect 281 74 285 78
rect -36 18 -32 22
rect 3 20 7 24
rect -10 13 -6 17
rect 23 13 27 17
rect 61 20 65 24
rect 49 13 53 17
rect 132 21 136 25
rect 171 20 175 24
rect 158 13 162 17
rect 191 13 195 17
rect 229 20 233 24
rect 217 13 221 17
rect 296 15 300 19
rect -86 -15 -82 -11
rect -68 -15 -64 -11
rect -52 -15 -48 -11
rect -28 -22 -24 -18
rect 99 -15 103 -11
rect 115 -15 119 -11
rect 40 -22 44 -18
rect 140 -22 144 -18
rect -18 -29 -14 -25
rect 31 -29 35 -25
rect 273 -15 277 -11
rect 209 -22 213 -18
rect 150 -29 154 -25
rect 199 -29 203 -25
<< ndcontact >>
rect -97 0 -93 4
rect -89 8 -85 12
rect -81 0 -77 4
rect -73 8 -69 12
rect -73 1 -69 5
rect -65 8 -61 12
rect -57 1 -53 5
rect -49 8 -45 12
rect -39 1 -35 5
rect -23 8 -19 12
rect 10 6 14 10
rect -7 1 -3 5
rect 20 1 24 5
rect 36 8 40 12
rect 68 6 72 10
rect 52 1 56 5
rect 96 0 100 4
rect 104 2 108 6
rect 112 8 116 12
rect 120 2 124 6
rect 129 1 133 5
rect 145 8 149 12
rect 178 6 182 10
rect 161 1 165 5
rect 188 1 192 5
rect 204 8 208 12
rect 236 6 240 10
rect 262 6 266 10
rect 270 8 274 12
rect 278 6 282 10
rect 286 8 290 12
rect 294 6 298 10
rect 302 8 306 12
rect 220 1 224 5
<< pdcontact >>
rect -97 59 -93 63
rect -73 27 -69 31
rect -49 59 -45 63
rect -39 45 -35 49
rect -23 29 -19 33
rect -7 45 -3 49
rect 20 45 24 49
rect 10 27 14 31
rect 36 29 40 33
rect 52 45 56 49
rect 78 39 82 43
rect 68 27 72 31
rect 86 45 90 49
rect 96 35 100 39
rect 104 27 108 31
rect 120 47 124 51
rect 129 45 133 49
rect 145 29 149 33
rect 161 45 165 49
rect 188 45 192 49
rect 178 27 182 31
rect 204 29 208 33
rect 262 59 266 63
rect 220 45 224 49
rect 246 39 250 43
rect 236 27 240 31
rect 254 45 258 49
rect 286 27 290 31
rect 294 35 298 39
rect 302 27 306 31
<< psubstratepcontact >>
rect -97 -8 -93 -4
rect -81 -8 -77 -4
rect -39 -8 -35 -4
rect -7 -8 -3 -4
rect 20 -8 24 -4
rect 52 -8 56 -4
rect 96 -8 100 -4
rect 129 -8 133 -4
rect 161 -8 165 -4
rect 188 -8 192 -4
rect 220 -8 224 -4
rect 262 -8 266 -4
rect 294 -8 298 -4
<< nsubstratencontact >>
rect -97 67 -93 71
rect -49 67 -45 71
rect -39 67 -35 71
rect 20 67 24 71
rect 86 67 90 71
rect 96 67 100 71
rect 120 67 124 71
rect 129 67 133 71
rect 188 67 192 71
rect 254 67 258 71
rect 262 67 266 71
rect 294 67 298 71
<< labels >>
rlabel metal1 -87 69 -87 69 5 vdd!
rlabel metal1 -98 74 -98 78 4 x
rlabel metal1 -82 74 -82 78 5 q0bar
rlabel metal1 -66 74 -66 78 5 q0
rlabel metal1 -87 -6 -87 -6 1 gnd!
rlabel metal1 -89 -15 -89 -11 1 q1
rlabel metal1 -43 18 -43 22 7 d0
rlabel metal1 -61 -15 -61 -11 1 q1bar
rlabel metal1 -45 -15 -45 -11 7 x
rlabel nsubstratencontact 98 69 98 69 4 vdd!
rlabel metal1 105 74 105 78 5 q0bar
rlabel psubstratepcontact 98 -6 98 -6 2 gnd!
rlabel metal1 97 -15 97 -11 2 xbar
rlabel metal1 113 -15 113 -11 1 q1
rlabel metal1 57 22 57 22 1 q0bar
rlabel metal1 78 16 78 20 1 q0
rlabel metal1 -29 -6 -29 -6 1 gnd!
rlabel metal1 -27 69 -27 69 1 vdd!
rlabel metal1 78 74 78 78 5 rst
rlabel metal1 139 -6 139 -6 1 gnd!
rlabel metal1 141 69 141 69 1 vdd!
rlabel metal1 246 74 246 78 5 rst
rlabel metal1 126 21 126 25 1 d1
rlabel metal1 246 16 246 20 1 q1
rlabel metal1 225 22 225 22 1 q1bar
rlabel metal1 277 74 277 78 5 q0bar
rlabel metal1 262 74 262 78 4 xbar
rlabel nsubstratencontact 264 69 264 69 4 vdd!
rlabel metal1 292 20 292 24 7 y
rlabel metal1 270 -15 270 -11 1 q1bar
rlabel psubstratepcontact 264 -6 264 -6 2 gnd!
rlabel metal1 295 15 295 19 1 x
rlabel metal1 308 15 308 19 7 xbar
rlabel metal1 -11 83 -11 83 1 clkbar
rlabel metal1 -17 90 -17 90 5 clk
<< end >>
